// Module:  complex_nr_mult_tb
// Author:  Gheorghe Stefan
// Date:    06.03.2020

module complex_nr_mult_tb(
    
);

endmodule // complex_nr_mult_tb