// Module:  clock_rst_gen
// Author:  Gheorghe Stefan
// Date:    06.03.2020

module clock_rst_gen(
    
);

endmodule // clock_rst_gen