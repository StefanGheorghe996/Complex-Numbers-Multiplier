//  Module: uint8_mult
//
module uint8_mult
    (
        input   [8 -1:0] op1,
        input   [8 -1:0] op2,
        output  [16-1:0] result
    );

    assign result =  op1 * op2;

    
endmodule
